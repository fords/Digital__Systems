library verilog;
use verilog.vl_types.all;
entity zxw_mux2to1_vlg_vec_tst is
end zxw_mux2to1_vlg_vec_tst;
