library verilog;
use verilog.vl_types.all;
entity zeyarW_lab1_vlg_vec_tst is
end zeyarW_lab1_vlg_vec_tst;
